module INV(
    output O,
    input I
);
  assign O = !I;
endmodule
